../../src_SSITH_P2/src_BSV/JtagTap.bsv