../../src_SSITH_P2/src_BSV/Giraffe_IFC.bsv