// Copyright (c) 2016-2021 Bluespec, Inc. All Rights Reserved.

// Widths of AXI buses

package AXI_Widths;

// ================================================================
// 'coherent DMA' port into L2 cache

typedef 16   Wd_Id_Dma;
typedef 64   Wd_Addr_Dma;
typedef 512  Wd_Data_Dma;
typedef 0    Wd_User_Dma;

// ================================================================

endpackage
