// Copyright (c) 2007--2011 Bluespec, Inc.  All rights reserved.
// $Revision$
// $Date$

package Axi;

////////////////////////////////////////////////////////////////////////////////
///
////////////////////////////////////////////////////////////////////////////////

import AxiDefines::*;
import AxiExtend::*;
import AxiMaster::*;
import AxiSlave::*;
import AxiRdBus::*;
import AxiWrBus::*;
import AxiPC::*;
// import AxiMonitor::*;

////////////////////////////////////////////////////////////////////////////////
///
////////////////////////////////////////////////////////////////////////////////

export AxiDefines::*;
export AxiExtend::*;
export AxiMaster::*;
export AxiSlave::*;
export AxiRdBus::*;
export AxiWrBus::*;
export AxiPC::*;
// export AxiMonitor::*;

endpackage
