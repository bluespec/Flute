../../src_SSITH_P2/src_BSV/ClockHacks.bsv